/////////////////////////////////////////////////////////////////                                               //
//    RISC-V                                                   //
//    RV12 Definitions Package                                 //
/////////////////////////////////////////////////////////////////

package riscv_rv12_pkg;
  parameter ARCHID       = 12;
  parameter REVPRV_MAJOR = 1;
  parameter REVPRV_MINOR = 10;
  parameter REVUSR_MAJOR = 2;
  parameter REVUSR_MINOR = 2;
endpackage

